
module esp 
#(
	parameter   clk_freq         = 100000000,
	parameter   uart_baud_rate   = 115200
)

(
	input CH_PD;
	input rx;
	output tx;
	input rst;

)





endmodule